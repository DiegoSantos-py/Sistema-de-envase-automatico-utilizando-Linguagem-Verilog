module MEF_main(
		input start, 
		input garrafa, 
		input sensor_de_nivel,
		input sensor_cq,
		input descarte,
		input ve_done,
		input cont_done,
		input clk,
		input reset,
		input alarme,
		output motor, 
		output EV,
		output pos_ve, // garrafa em posição de vedação
		output count, // sinal para ativar mef do contador
		output resetar,
		output Desc_signal,
		output controle_qualidade,
		output pos_cq
		);
		
		reg[2:0]state, nextstate;
		
		parameter SR = 3'b000; // Start/reset
		parameter Mo = 3'b001; // Motor
		parameter En = 3'b010; // Enchimento
		parameter Vd = 3'b011; // Vedação
		parameter Cq = 3'b100; // Controle de qualidade
		parameter Co = 3'b101; // Contador
		parameter De = 3'b110; // Descarte
		
		always @ ( posedge clk , posedge
		reset )
			if ( reset ) state <= SR ;
			else state <= nextstate ;
			
		always @(*)
			case(state)
				SR:
					nextstate = Mo;
				Mo:
					if (start == 1)
						nextstate = SR;
					else if (alarme == 1)
						nextstate = Mo;
					else if (garrafa == 1)
						nextstate = En;
					else
						nextstate = Mo;
				En:
					if (start == 1)
						nextstate = SR;
					else if (sensor_de_nivel == 1) 
						nextstate = Vd;
					else
						nextstate = En;
				Vd:
					if (start == 1)
						nextstate = SR;
					else if (ve_done == 1)
						nextstate = Cq;
					else
						nextstate = Vd;
				Cq:
					if (start == 1)
						nextstate = SR;
					else if (sensor_cq == 1)
						nextstate = Co;
					else if (descarte == 1)
						nextstate = De;
					else
						nextstate = Cq;
				Co:
					if (start == 1)
						nextstate = SR;
					else if (cont_done == 1)
						nextstate = Mo;
					else
						nextstate = Co;
				De:
					nextstate = Mo;
				default:
                nextstate = SR;
			endcase
		
		// Motor deve ficar ligado quando tiver garrafa e mef está em Mo
		assign resetar = (state == SR);
		assign motor = (state == Mo);
		assign EV = (state == En);
		assign pos_ve = (state == Vd);
		assign controle_qualidade = (state == Cq);
		assign count = (state == Co);
		assign Desc_signal = (state == De);
		assign pos_cq = (state == Cq);

endmodule