module d_flipflop (
    input d,
    input  clk,
    input  reset,
    output wire q
);
	wire nreset;
	not(nreset, reset);
	dff flipflop_inst (
		 .d(d),
		 .clk(clk),
		 .clrn(nreset),  
		 .q(q)
);

endmodule